//@author christian yu 104785497
`include "led_fsm.v"
`include "code_reg.v"
////////////////////////////////////////////////////////////////
//  Main File for dassign3 
////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////
//  module dassign3 (also MORSE_ENCODER)
////////////////////////////////////////////////////////////////
module dassign3(
		input 	    char_vald,
		input [7:0] charcode_data,
		input [3:0] charlen_data,
		output 	    char_next, led_drv,
		input 	    reset, clock
		);

////////////////////////////////////////////////////////////////
//  Parameter Declarations
////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////
//  Variable Declaration
////////////////////////////////////////////////////////////////

   // Outputs from modules       
   wire       shft_data, sym_done, led_drv; 
   wire [3:0] cntr_data; 

   // Signals that needs to be generated by this module
   reg 	      char_next, char_load, shft_cnt, sym_strt;

////////////////////////////////////////////////////////////////
//  Module Instantiation
////////////////////////////////////////////////////////////////

   code_reg codestore0(charcode_data, charlen_data, char_load, 
                       sym_done, cntr_data, shft_data, reset, clock);
   led_fsm ledfsm0(sym_strt, shft_data, led_drv, sym_done, 
                   reset, clock);
        
/* Some useful pseudo-code (you have to figure out if there are
   timing consideration or sequencing that you would want to do.
   From that, you can choose to build an FSM. You can choose to 
   build it as a separate module).
 
 symbol for led_fsm = shft_data from the shifter
 sym_strt is asserted when char_vald or after you've shifted 
    a new data symbol from the shifter

 space symbol is detected when charlen_data = 4'b0000      
 shft_cnt is asserted when sym_done is asserted (if using the 
    counter to deal with a space, you'd need to enable shft_cnt for 
    a "space" symbol)

 char_next for encoder = cntr counts down to 0
    (load counter with 4'b0111 when it is a space either in 
    code_reg or here)
 char_ vald input should trigger the char_load to grab the new 
    charcode_data and charlen_data
 */

////////////////////////////////////////////////////////////////
//  STATE MACHINE
////////////////////////////////////////////////////////////////
  
  reg [3:0] morse_st, morse_nx_st;
  
  parameter IDLE = 4'b0000;
  parameter LOAD = 4'b0001;
  parameter CHAR = 4'b0011;
  parameter BLNK1= 4'b0010;
  parameter BLNK2= 4'b0110;
  parameter BLNK3= 4'b0111;
  parameter BLNK4= 4'b0101;
  parameter BLNK5= 4'b0100;
  parameter BLNK6= 4'b1100;
  parameter BLNK7= 4'b1000;
  
  always @(posedge clock) begin
    morse_st <= morse_nx_st;
  end
  
////////////////////////////////////////////////////////////////
//  FSM LOGIC
////////////////////////////////////////////////////////////////  
  
  always @(*) begin
    if(reset) begin
      morse_nx_st = IDLE;
      char_next = 1;
      char_load = 0;
      sym_strt  = 0;
    end
    
    else begin
      case(morse_st)
        IDLE: begin
          if(char_vald) begin
            char_next = 0;
            if(charlen_data == 4'b0000) begin
              char_load = 0;
              morse_nx_st = BLNK1;
            end
            else begin
              char_load = 1;
              morse_nx_st = LOAD;
            end
          end
          else begin
            morse_nx_st = IDLE;
            char_next = 1;
            char_load = 0;
          end
        end
        
        LOAD: begin
            char_load = 0;
            morse_nx_st = CHAR;
        end
        
        CHAR: begin
          if(cntr_data == 4'b0000) begin
          	sym_strt = 0;
            morse_nx_st = IDLE;
            char_next = 1;
          end
          else begin
            sym_strt = 1;
            morse_nx_st = CHAR;
          end
        end
        
        BLNK1: begin
          morse_nx_st = BLNK2;
        end
        BLNK2: begin
          morse_nx_st = BLNK3;
        end
        BLNK3: begin
          morse_nx_st = BLNK4;
        end
        BLNK4: begin
          morse_nx_st = BLNK5;
        end
        BLNK5: begin
          morse_nx_st = BLNK6;
        end
        BLNK6: begin
          morse_nx_st = BLNK7;
        end
        BLNK7: begin
          morse_nx_st = IDLE;
          char_next = 1;
        end
        
        default: begin
     	 morse_nx_st = IDLE;
     	 char_next = 1;
    	 char_load = 0;
     	 sym_strt  = 0;
        end
      endcase
    end
  end
    
endmodule // dassign3